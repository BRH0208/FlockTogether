{"tileData":"{\"seed\":2658,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":40.75188064575195,\"y\":34.68705368041992},{\"x\":40.214542388916019,\"y\":34.59286880493164},{\"x\":40.26117706298828,\"y\":34.3875846862793},{\"x\":40.72446823120117,\"y\":34.95371627807617},{\"x\":40.33146286010742,\"y\":34.25631332397461},{\"x\":40.75188064575195,\"y\":34.68705368041992},{\"x\":40.214542388916019,\"y\":34.59286880493164},{\"x\":40.26117706298828,\"y\":34.3875846862793},{\"x\":40.72446823120117,\"y\":34.95371627807617},{\"x\":40.33146286010742,\"y\":34.25631332397461}]}"],"dataNames":["ZMan"]}