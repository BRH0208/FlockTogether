{"tileData":"{\"seed\":3035,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":37.435203552246097,\"y\":39.24506378173828},{\"x\":37.79424285888672,\"y\":39.592185974121097},{\"x\":37.63746643066406,\"y\":39.16842269897461},{\"x\":37.75040817260742,\"y\":39.697242736816409},{\"x\":37.03464126586914,\"y\":39.93101119995117},{\"x\":37.435203552246097,\"y\":39.24506378173828},{\"x\":37.79424285888672,\"y\":39.592185974121097},{\"x\":37.63746643066406,\"y\":39.16842269897461},{\"x\":37.75040817260742,\"y\":39.697242736816409},{\"x\":37.03464126586914,\"y\":39.93101119995117}]}"],"dataNames":["ZMan"]}