{"tileData":"{\"seed\":2656,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":38.128814697265628,\"y\":34.83610534667969},{\"x\":38.37287139892578,\"y\":34.48055648803711},{\"x\":38.38837814331055,\"y\":34.565338134765628},{\"x\":38.128814697265628,\"y\":34.83610534667969},{\"x\":39.10592269897461,\"y\":34.64132308959961},{\"x\":38.00102233886719,\"y\":35.064781188964847},{\"x\":38.37287139892578,\"y\":34.48055648803711},{\"x\":38.38837814331055,\"y\":34.565338134765628}]}"],"dataNames":["ZMan"]}