{"tileData":"{\"seed\":2655,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":37.5512580871582,\"y\":34.3894157409668},{\"x\":37.23515319824219,\"y\":34.10823059082031},{\"x\":37.332191467285159,\"y\":34.939884185791019},{\"x\":37.28449630737305,\"y\":34.60627365112305},{\"x\":37.47537612915039,\"y\":34.041927337646487},{\"x\":37.5512580871582,\"y\":34.3894157409668},{\"x\":37.23515319824219,\"y\":34.10823059082031},{\"x\":37.332191467285159,\"y\":34.939884185791019},{\"x\":37.28449630737305,\"y\":34.60627365112305},{\"x\":37.47537612915039,\"y\":34.041927337646487},{\"x\":37.62502670288086,\"y\":34.9014892578125},{\"x\":37.868316650390628,\"y\":34.88175964355469}]}"],"dataNames":["ZMan"]}