{"tileData":"{\"seed\":2581,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":39.834327697753909,\"y\":33.835044860839847},{\"x\":39.08436584472656,\"y\":33.333248138427737},{\"x\":39.41682815551758,\"y\":33.165794372558597},{\"x\":39.65913772583008,\"y\":33.29964828491211},{\"x\":39.413909912109378,\"y\":33.61717987060547},{\"x\":39.834327697753909,\"y\":33.835044860839847},{\"x\":39.08436584472656,\"y\":33.333248138427737},{\"x\":39.41682815551758,\"y\":33.165794372558597},{\"x\":39.65913772583008,\"y\":33.29964828491211},{\"x\":39.413909912109378,\"y\":33.61717987060547}]}"],"dataNames":["ZMan"]}