{"tileData":"{\"seed\":2580,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":38.6715202331543,\"y\":33.63236618041992},{\"x\":38.48931884765625,\"y\":33.4792594909668},{\"x\":38.551429748535159,\"y\":33.19093322753906},{\"x\":38.947998046875,\"y\":33.58531188964844},{\"x\":38.21336364746094,\"y\":33.750205993652347},{\"x\":38.6715202331543,\"y\":33.63236618041992},{\"x\":38.48931884765625,\"y\":33.4792594909668},{\"x\":38.551429748535159,\"y\":33.19093322753906},{\"x\":38.947998046875,\"y\":33.58531188964844},{\"x\":38.21336364746094,\"y\":33.750205993652347}]}"],"dataNames":["ZMan"]}