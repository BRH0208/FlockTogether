{"tileData":"{\"seed\":3037,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":39.108123779296878,\"y\":39.3618049621582},{\"x\":39.9885368347168,\"y\":39.89120864868164},{\"x\":39.80046844482422,\"y\":39.762428283691409},{\"x\":39.048038482666019,\"y\":39.56110763549805},{\"x\":39.070899963378909,\"y\":39.719024658203128},{\"x\":39.108123779296878,\"y\":39.3618049621582},{\"x\":39.9885368347168,\"y\":39.89120864868164},{\"x\":39.80046844482422,\"y\":39.762428283691409},{\"x\":39.048038482666019,\"y\":39.56110763549805},{\"x\":39.070899963378909,\"y\":39.719024658203128}]}"],"dataNames":["ZMan"]}