{"tileData":"{\"seed\":2730,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":36.9238395690918,\"y\":35.25674057006836},{\"x\":36.71999740600586,\"y\":35.96662521362305},{\"x\":36.22147750854492,\"y\":35.21523666381836},{\"x\":36.83387756347656,\"y\":35.364654541015628},{\"x\":36.826290130615237,\"y\":35.50291061401367},{\"x\":36.9238395690918,\"y\":35.25674057006836},{\"x\":36.71999740600586,\"y\":35.96662521362305},{\"x\":36.22147750854492,\"y\":35.21523666381836},{\"x\":36.83387756347656,\"y\":35.364654541015628},{\"x\":36.826290130615237,\"y\":35.50291061401367}]}"],"dataNames":["ZMan"]}