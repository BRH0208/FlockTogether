{"tileData":"{\"seed\":3036,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":38.50725555419922,\"y\":39.60836410522461},{\"x\":38.59947967529297,\"y\":39.09020233154297},{\"x\":38.72734069824219,\"y\":39.871009826660159},{\"x\":38.526954650878909,\"y\":39.58274459838867},{\"x\":38.628421783447269,\"y\":39.42182540893555},{\"x\":38.50725555419922,\"y\":39.60836410522461},{\"x\":38.59947967529297,\"y\":39.09020233154297},{\"x\":38.72734069824219,\"y\":39.871009826660159},{\"x\":38.526954650878909,\"y\":39.58274459838867},{\"x\":38.628421783447269,\"y\":39.42182540893555}]}"],"dataNames":["ZMan"]}