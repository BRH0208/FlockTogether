{"tileData":"{\"seed\":3112,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":38.02569580078125,\"y\":40.57132339477539},{\"x\":38.779632568359378,\"y\":40.372989654541019},{\"x\":38.4054069519043,\"y\":40.666751861572269},{\"x\":38.66828155517578,\"y\":40.97394561767578},{\"x\":38.23739242553711,\"y\":40.15195083618164},{\"x\":38.02569580078125,\"y\":40.57132339477539},{\"x\":38.779632568359378,\"y\":40.372989654541019},{\"x\":38.4054069519043,\"y\":40.666751861572269},{\"x\":38.66828155517578,\"y\":40.97394561767578},{\"x\":38.23739242553711,\"y\":40.15195083618164}]}"],"dataNames":["ZMan"]}