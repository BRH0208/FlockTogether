{"tileData":"{\"seed\":2657,\"didGenerate\":true}","data":["{\"zombies\":[{\"x\":39.387359619140628,\"y\":34.918216705322269},{\"x\":39.32130432128906,\"y\":34.03450393676758},{\"x\":39.699466705322269,\"y\":34.10227966308594},{\"x\":39.713584899902347,\"y\":34.82394790649414},{\"x\":39.44106674194336,\"y\":34.99993896484375},{\"x\":39.387359619140628,\"y\":34.918216705322269},{\"x\":39.32130432128906,\"y\":34.03450393676758},{\"x\":39.699466705322269,\"y\":34.10227966308594},{\"x\":39.713584899902347,\"y\":34.82394790649414},{\"x\":39.75883865356445,\"y\":34.97721481323242},{\"x\":39.411651611328128,\"y\":34.79022979736328},{\"x\":39.10592269897461,\"y\":34.64132308959961},{\"x\":39.44106674194336,\"y\":34.99993896484375}]}"],"dataNames":["ZMan"]}